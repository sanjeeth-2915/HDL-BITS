module top_module( 
    input a,b,c,
    output w,x,y,z );
	//initial begin 
      assign w=a; 
      assign x=b,y=b; 
        
       assign z=c;
   // end
endmodule
